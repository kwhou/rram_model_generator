.subckt cell TE BE RM=10K
* X1  TE   BE   rram
R1  TE   BE   'RM'
.ends
